module latch_8bit (
    input               rst_n,
    input [7:0]         data_8b_in,
    input               data_en,
    output reg [7:0]    data_8b_out
);
    reg [7:0]          bus_net0;

    always @ (*) begin
        if (!rst_n) begin
            data_8b_out = 8'h00;
            bus_net0    = 8'h00;
        end
        else begin
            if (data_en) begin
                data_8b_out = data_8b_in;
                bus_net0    = 8'h00;
            end
            else begin
                bus_net0    = data_8b_out;
                data_8b_out = bus_net0;
            end
        end
    end

endmodule